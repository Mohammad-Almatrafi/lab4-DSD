`timescale 1ns / 1ps

module mult_8bit(

    );
endmodule
